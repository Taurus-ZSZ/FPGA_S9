module S9_top(


);



endmodule
